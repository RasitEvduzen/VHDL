exp1_inst : exp1 PORT MAP (
		aclr	 => aclr_sig,
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
